`timescale 1ns/1ps




module RegisterFile(A1,A2,A3,WD3,clk, WE3,RD1, RD2, rst, RD3); // A3 is the destination regiter.
    input [4:0] A1,A2,A3;
    input [31:0]WD3;
    input clk, WE3, rst;
    output [31:0] RD1, RD2, RD3;
    
    integer i;
    reg [31:0] mem[0:31];
    reg [31:0] mem_next;
    
    assign RD3 = mem[7];
    
//    initial begin
//        $readmemh("reg_mem.mem", mem);
//        end
    always @(negedge clk )begin
        if (WE3 == 1 && A3 != 32'b0)     // Because register zero is only to store zero values.                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          
            mem[A3] <= WD3;
        else 
            mem[A3] <= mem_next;
    end
    
    // Hold the prvous state.
    always@ (*) begin
        mem_next = mem[A3];
    end 
    
    assign RD1 = rst? 32'b0 : mem[A1];
    assign RD2 = rst? 32'b0 : mem[A2];
    
    initial begin
        mem[0] = 32'b0;
        mem[1] = 32'h5;
        mem[5] = 32'h6;
        mem[7] = 32'h9;
        mem[6] = 32'ha;
        mem[4] = 32'h1;
        mem[19] = 32'b1;
        mem[20] = 32'h4;
        mem[8] = 32'h456;
        mem[9] = 32'h2004;
        mem[21] = 32'h0;
        mem[28] = 32'h9;
       end
endmodule
